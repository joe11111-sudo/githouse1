library verilog;
use verilog.vl_types.all;
entity mips is
end mips;
